
module decoder5to32(enable, select, out_add);
    input           enable;
    input   [4:0]   select;
    output reg [31:0]  out_add;
 
always @(*) 
    begin
    if (enable) 
        begin
            case(select)
                5'b00000: out_add = 32'b0000_0000_0000_0000_0000_0000_0000_0001;
                5'b00001: out_add = 32'b0000_0000_0000_0000_0000_0000_0000_0010;
                5'b00010: out_add = 32'b0000_0000_0000_0000_0000_0000_0000_0100;
                5'b00011: out_add = 32'b0000_0000_0000_0000_0000_0000_0000_1000;
                5'b00100: out_add = 32'b0000_0000_0000_0000_0000_0000_0001_0000;
                5'b00101: out_add = 32'b0000_0000_0000_0000_0000_0000_0010_0000;
                5'b00110: out_add = 32'b0000_0000_0000_0000_0000_0000_0100_0000;
                5'b00111: out_add = 32'b0000_0000_0000_0000_0000_0000_1000_0000;
                5'b01000: out_add = 32'b0000_0000_0000_0000_0000_0001_0000_0000;
                5'b01001: out_add = 32'b0000_0000_0000_0000_0000_0010_0000_0000;
                5'b01010: out_add = 32'b0000_0000_0000_0000_0000_0100_0000_0000;
                5'b01011: out_add = 32'b0000_0000_0000_0000_0000_1000_0000_0000;
                5'b01100: out_add = 32'b0000_0000_0000_0000_0001_0000_0000_0000;
                5'b01101: out_add = 32'b0000_0000_0000_0000_0010_0000_0000_0000;
                5'b01110: out_add = 32'b0000_0000_0000_0000_0100_0000_0000_0000;
                5'b01111: out_add = 32'b0000_0000_0000_0000_1000_0000_0000_0000;
                
                5'b10000: out_add = 32'b0000_0000_0000_0001_0000_0000_0000_0000;
                5'b10001: out_add = 32'b0000_0000_0000_0010_0000_0000_0000_0000;
                5'b10010: out_add = 32'b0000_0000_0000_0100_0000_0000_0000_0000;
                5'b10011: out_add = 32'b0000_0000_0000_1000_0000_0000_0000_0000;
                5'b10100: out_add = 32'b0000_0000_0001_0000_0000_0000_0000_0000;
                5'b10101: out_add = 32'b0000_0000_0010_0000_0000_0000_0000_0000;
                5'b10110: out_add = 32'b0000_0000_0100_0000_0000_0000_0000_0000;
                5'b10111: out_add = 32'b0000_0000_1000_0000_0000_0000_0000_0000;
                5'b11000: out_add = 32'b0000_0001_0000_0000_0000_0000_0000_0000;
                5'b11001: out_add = 32'b0000_0010_0000_0000_0000_0000_0000_0000;
                5'b11010: out_add = 32'b0000_0100_0000_0000_0000_0000_0000_0000;
                5'b11011: out_add = 32'b0000_1000_0000_0000_0000_0000_0000_0000;
                5'b11100: out_add = 32'b0001_0000_0000_0000_0000_0000_0000_0000;
                5'b11101: out_add = 32'b0010_0000_0000_0000_0000_0000_0000_0000;
                5'b11110: out_add = 32'b0100_0000_0000_0000_0000_0000_0000_0000;
                5'b11111: out_add = 32'b1000_0000_0000_0000_0000_0000_0000_0000;
            endcase
        end
    else
        out_add = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    end

endmodule