module OR_Gate(A, B, O);
input A, B;
output O

assign 0 = A | B;

endmodule